library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VGA_green is
	port(	CLOCK_50 : in std_logic; -- clock interne
			KEY     : in std_logic_vector(3 downto 0); -- bouton
			SW      : in std_logic_vector(9 downto 0); -- switch
			VGA_R, VGA_G, VGA_B : out std_logic_vector(3 downto 0); -- signaux RGB du ADV7123
			VGA_CLK : inout std_logic;  -- signaux du MAX10
			BLANK_N : out std_logic;-- signaux du MAX10
			VGA_HS  : out std_logic;-- signaux du MAX10
			VGA_VS  : out std_logic;-- signaux du MAX10
			GPIO    : out std_logic_vector(34 downto 0)
	);
end entity;

architecture DE1_SoC of VGA_green is
	
	component pll_vga is
		port 	(
			inclk0	: IN STD_LOGIC  := '0';
			c0		   : OUT STD_LOGIC 
		);
	end component pll_vga;	

	signal reset : std_logic;

begin

----------------------------------------------------------------
-- port map du pll
----------------------------------------------------------------
	
	pll : pll_vga port map (
		inclk0 => CLOCK_50,
		c0		 => VGA_CLK
	);
	
----------------------------------------------------------------
-- Définir la couleur
----------------------------------------------------------------

	reset <= not KEY(0);

	GPIO(0) <= VGA_CLK;
	
----------------------------------------------------------------
-- Générer les signaux de sync
----------------------------------------------------------------
   process(VGA_CLK, KEY(0)) is
      variable hcount : integer range 0 to 800;
      variable vcount : integer range 0 to 525;
   begin
	
		-- RESET
      if(KEY(0) = '0') then
         hcount := 0;
         vcount := 0;
         vga_hs <= '1';
         vga_vs <= '1';
			BLANK_N  <= '0';
			
      elsif(VGA_CLK'event and VGA_CLK = '1') then

         if(hcount >= 0 and hcount <= 639 and vcount >= 0 and vcount <= 479) then
				VGA_R <= "1111";
				VGA_G <= "0000";
				VGA_B <= "0000";
		
         else
			-- blank the screen when not in range
				VGA_R <= "0000";
				VGA_G <= "0000";
				VGA_B <= "0000";

			end if;
			
			-- Incrémente les compteurs hcount / vcount
			if(hcount = 799) then
				hcount := 0;
				if(vcount = 524) then	
					vcount := 0;
				else
					vcount := vcount + 1;
				end if;
			else
				hcount := hcount + 1;
			end if;
			
			-- Définit le sync pulse horizontal
			if(hcount = 656) then		vga_hs <= '0';
			elsif(hcount = 752) then	vga_hs <= '1';
			end if;
			
			-- Définit le sync pulse vertical
			if(vcount = 490) then		vga_vs <= '0';
			elsif(vcount = 492) then	vga_vs <= '1';
			end if;
			
      end if;
   end process;
	
end DE1_SoC;
